*** multiStage.cir ***
* Shared nodes:  gnd, cc (+12V), ee (-12V), s, in, out
* Stage 1 nodes: e1, c1
* Stage 2 nodes: b2, e2, e22, c2
* Stage 3 nodes: b3, e3, e33, c3
* Stage 4 nodes: b4, e4
*
*POWER SUPPLIES AND SOURCE
Vcc cc gnd dc 12V ac 0V
Vee ee gnd dc -12V ac 0V
Vs s gnd dc 0V ac 10mV
Rs in s 50
*
*STAGE 1; COMMON BASE
Cc1 in e1 3.183uF
Re1 e1 ee 21.8k
Q1 c1 gnd e1 model1
L1 c1 cc 3.0uH
Cd1 c1 cc 80pF
Rp1 c1 cc 21.7k 
*
*STAGE 2: COMMON EMITTER
Cc2 c1 b2 11.4nF
R1 cc b2 378.9k
R2 b2 ee 425.8k
Q2 c2 b2 e2 model2
Rex2 e2 e22 50
Re2 e22 ee 10.5k
Ce2 e22 gnd 25.5nF
L2 c2 cc 4.2uH
Cd2 c2 cc 61.66pF
Rp2 c2 cc 40.3k
*
*STAGE 3: COMMON EMITTER
Cc3 c2 b3 11.4nF
R3 cc b3 378.9k
R4 b3 ee 425.8k
Q3 c3 b3 e3 model3
Rex3 e3 e33 50
Re3 e33 ee 10.5k
Ce3 e33 gnd 25.5nF
L3 c3 cc 4.4uH
Cd3 c3 cc 64.33pF
Rp3 c3 cc 30.4k
*
*STAGE 4: COMMON COLLECTOR
Cc4 c3 b4 13nF
R5 cc b4 833k
R6 b4 ee 936.2k
Q4 cc b4 e4 model4
Re4 e4 ee 23.2k
*
*OUTPUT
Cc5 e4 out 3.18iuF
Rload out gnd 100k
*
* .model <name> <type> (par1=value1 par2=value2 ...)
* VAF = forward Early voltage
* BF = forward beta; forward common-emitter gain
* CJE = base-emitter zero-bias junction capacitance
* CJC = base-collector zero-bias junction capacitance
* TS = transport saturation current
* NF = forward mode ideality factor
*
.model model1 npn (BF=181 CJC=5.1pf CJE=3.26pf IS=1E-16 VAF=260V NF=1)
.model model2 npn (BF=191 CJC=5.19pf CJE=3.28pf IS=1E-16 VAF=273V NF=1) ; CJC has large effect on CB gain and CC2 throughput
.model model3 npn (BF=189 CJC=5.18pf CJE=3.30pf IS=1E-16 VAF=273V NF=1)
.model model4 npn (BF=189 CJC=5.23pf CJE=3.24pf IS=1E-16 VAF=224V NF=1) ; model2 CJE has effect on CC2 throughput but not CB gain
*
*OUTPUT CONTROL
.control
set filetype=ascii
.op
*ac dec 10 1Hz 1GHz
ac dec 10 100kHz 1GHz
plot db(v(out)/v(in))
plot ph(v(out))-ph(v(in))
write multiStage.txt db(v(out)/v(in)) ph(v(out))-ph(v(in))

