*** CBstage.cir ***
* Nodes:
* gnd, cc (+12V), ee (-12V), s, in, e1, c1, out

Vcc cc gnd dc 12V ac 0V
Vee ee gnd dc -12V ac 0V
Vs s gnd dc 0V ac 10mV
Rs in s 50
Cc1 in e1 3.183uF
Re1 e1 ee 21.8k
Q1 c1 gnd e1 model1
L1 c1 cc 4.2uH
Cd1 c1 cc 55pF
Rp1 c1 cc 2.18k
Cc2 c1 out 3.183uF
Rld out gnd 9999k

* .model <name> <type> (par1=value1 par2=value2 ...)
* VAF = forward Early voltage
* BF = forward beta; forward common-emitter gain
* CJE = base-emitter zero-bias junction capacitance
* CJC = base-collector zero-bias junction capacitance
* TS = transport saturation current
* NF = forward mode ideality factor

.model model1 npn (BF=176 CJC=20pf CJE=20pf IS=1E-16 VAF=452V NF=1)

.control
set filetype=ascii
ac dec 10 1Hz 1GHz
plot db(v(out)/v(in))
plot ph(v(out))-ph(v(in))
write CBstage.txt db(v(output)/v(input)) ph(v(output))-ph(v(input))

