*** multiStage.cir ***
* Nodes:
* gnd, cc (+12V), ee (-12V), s, in, b2, e2, e22, c2, out

Vcc cc gnd dc 12V ac 0V
Vee ee gnd dc -12V ac 0V
Vs s gnd dc 0V ac 10mV
Rs in s 50
Cc2 in b2 13nF
R1 cc b2 177.2k
R2 b2 ee 96.6k
Q2 c2 b2 e2 model2
Rex e2 e22 50
Re2 e22 ee 6.25k
Ce2 e22 gnd 25.5nF
L2 c2 cc 4.2uH
Cd2 c2 cc 55pF
Rp2 c2 cc 30k
Cc3 c2 out 13nF
Rld out gnd 9999k

* .model <name> <type> (par1=value1 par2=value2 ...)
* VAF = forward Early voltage
* BF = forward beta; forward common-emitter gain
* CJE = base-emitter zero-bias junction capacitance
* CJC = base-collector zero-bias junction capacitance
* TS = transport saturation current
* NF = forward mode ideality factor

.model model2 npn (BF=192 CJC=20pf CJE=20pf IS=1E-16 VAF=228V NF=1)

.control
set filetype=ascii
ac dec 10 1Hz 1GHz
plot db(v(out)/v(s))
plot ph(v(out))-ph(v(s))
write CEstage.txt db(v(out)/v(s)) ph(v(out))-ph(v(s))

.end
